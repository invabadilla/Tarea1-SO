// platform.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module platform (
		input  wire        clk_clk,                                  //                               clk.clk
		output wire [13:0] id7segm_min_0_external_connection_export, // id7segm_min_0_external_connection.export
		output wire [13:0] id7segm_ms_0_external_connection_export,  //  id7segm_ms_0_external_connection.export
		output wire [13:0] id7segm_s_0_external_connection_export,   //   id7segm_s_0_external_connection.export
		input  wire [1:0]  pio_0_external_connection_export,         //         pio_0_external_connection.export
		input  wire        reset_reset_n,                            //                             reset.reset_n
		input  wire [2:0]  switches_0_external_connection_export     //    switches_0_external_connection.export
	);

	wire  [31:0] cpu_0_data_master_readdata;                 // mm_interconnect_0:CPU_0_data_master_readdata -> CPU_0:d_readdata
	wire         cpu_0_data_master_waitrequest;              // mm_interconnect_0:CPU_0_data_master_waitrequest -> CPU_0:d_waitrequest
	wire  [14:0] cpu_0_data_master_address;                  // CPU_0:d_address -> mm_interconnect_0:CPU_0_data_master_address
	wire   [3:0] cpu_0_data_master_byteenable;               // CPU_0:d_byteenable -> mm_interconnect_0:CPU_0_data_master_byteenable
	wire         cpu_0_data_master_read;                     // CPU_0:d_read -> mm_interconnect_0:CPU_0_data_master_read
	wire         cpu_0_data_master_write;                    // CPU_0:d_write -> mm_interconnect_0:CPU_0_data_master_write
	wire  [31:0] cpu_0_data_master_writedata;                // CPU_0:d_writedata -> mm_interconnect_0:CPU_0_data_master_writedata
	wire         mm_interconnect_0_ram_0_s1_chipselect;      // mm_interconnect_0:RAM_0_s1_chipselect -> RAM_0:chipselect
	wire  [31:0] mm_interconnect_0_ram_0_s1_readdata;        // RAM_0:readdata -> mm_interconnect_0:RAM_0_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_0_s1_address;         // mm_interconnect_0:RAM_0_s1_address -> RAM_0:address
	wire   [3:0] mm_interconnect_0_ram_0_s1_byteenable;      // mm_interconnect_0:RAM_0_s1_byteenable -> RAM_0:byteenable
	wire         mm_interconnect_0_ram_0_s1_write;           // mm_interconnect_0:RAM_0_s1_write -> RAM_0:write
	wire  [31:0] mm_interconnect_0_ram_0_s1_writedata;       // mm_interconnect_0:RAM_0_s1_writedata -> RAM_0:writedata
	wire         mm_interconnect_0_ram_0_s1_clken;           // mm_interconnect_0:RAM_0_s1_clken -> RAM_0:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;    // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;      // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;       // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;         // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;     // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] mm_interconnect_0_switches_0_s1_readdata;   // switches_0:readdata -> mm_interconnect_0:switches_0_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_0_s1_address;    // mm_interconnect_0:switches_0_s1_address -> switches_0:address
	wire         mm_interconnect_0_buttons_0_s1_chipselect;  // mm_interconnect_0:buttons_0_s1_chipselect -> buttons_0:chipselect
	wire  [31:0] mm_interconnect_0_buttons_0_s1_readdata;    // buttons_0:readdata -> mm_interconnect_0:buttons_0_s1_readdata
	wire   [1:0] mm_interconnect_0_buttons_0_s1_address;     // mm_interconnect_0:buttons_0_s1_address -> buttons_0:address
	wire         mm_interconnect_0_buttons_0_s1_write;       // mm_interconnect_0:buttons_0_s1_write -> buttons_0:write_n
	wire  [31:0] mm_interconnect_0_buttons_0_s1_writedata;   // mm_interconnect_0:buttons_0_s1_writedata -> buttons_0:writedata
	wire         mm_interconnect_0_segm_ms_0_s1_chipselect;  // mm_interconnect_0:segm_ms_0_s1_chipselect -> segm_ms_0:chipselect
	wire  [31:0] mm_interconnect_0_segm_ms_0_s1_readdata;    // segm_ms_0:readdata -> mm_interconnect_0:segm_ms_0_s1_readdata
	wire   [1:0] mm_interconnect_0_segm_ms_0_s1_address;     // mm_interconnect_0:segm_ms_0_s1_address -> segm_ms_0:address
	wire         mm_interconnect_0_segm_ms_0_s1_write;       // mm_interconnect_0:segm_ms_0_s1_write -> segm_ms_0:write_n
	wire  [31:0] mm_interconnect_0_segm_ms_0_s1_writedata;   // mm_interconnect_0:segm_ms_0_s1_writedata -> segm_ms_0:writedata
	wire         mm_interconnect_0_segm_s_0_s1_chipselect;   // mm_interconnect_0:segm_s_0_s1_chipselect -> segm_s_0:chipselect
	wire  [31:0] mm_interconnect_0_segm_s_0_s1_readdata;     // segm_s_0:readdata -> mm_interconnect_0:segm_s_0_s1_readdata
	wire   [1:0] mm_interconnect_0_segm_s_0_s1_address;      // mm_interconnect_0:segm_s_0_s1_address -> segm_s_0:address
	wire         mm_interconnect_0_segm_s_0_s1_write;        // mm_interconnect_0:segm_s_0_s1_write -> segm_s_0:write_n
	wire  [31:0] mm_interconnect_0_segm_s_0_s1_writedata;    // mm_interconnect_0:segm_s_0_s1_writedata -> segm_s_0:writedata
	wire         mm_interconnect_0_segm_min_0_s1_chipselect; // mm_interconnect_0:segm_min_0_s1_chipselect -> segm_min_0:chipselect
	wire  [31:0] mm_interconnect_0_segm_min_0_s1_readdata;   // segm_min_0:readdata -> mm_interconnect_0:segm_min_0_s1_readdata
	wire   [1:0] mm_interconnect_0_segm_min_0_s1_address;    // mm_interconnect_0:segm_min_0_s1_address -> segm_min_0:address
	wire         mm_interconnect_0_segm_min_0_s1_write;      // mm_interconnect_0:segm_min_0_s1_write -> segm_min_0:write_n
	wire  [31:0] mm_interconnect_0_segm_min_0_s1_writedata;  // mm_interconnect_0:segm_min_0_s1_writedata -> segm_min_0:writedata
	wire  [31:0] cpu_0_instruction_master_readdata;          // mm_interconnect_1:CPU_0_instruction_master_readdata -> CPU_0:i_readdata
	wire         cpu_0_instruction_master_waitrequest;       // mm_interconnect_1:CPU_0_instruction_master_waitrequest -> CPU_0:i_waitrequest
	wire  [14:0] cpu_0_instruction_master_address;           // CPU_0:i_address -> mm_interconnect_1:CPU_0_instruction_master_address
	wire         cpu_0_instruction_master_read;              // CPU_0:i_read -> mm_interconnect_1:CPU_0_instruction_master_read
	wire         mm_interconnect_1_rom_0_s1_chipselect;      // mm_interconnect_1:ROM_0_s1_chipselect -> ROM_0:chipselect
	wire  [31:0] mm_interconnect_1_rom_0_s1_readdata;        // ROM_0:readdata -> mm_interconnect_1:ROM_0_s1_readdata
	wire         mm_interconnect_1_rom_0_s1_debugaccess;     // mm_interconnect_1:ROM_0_s1_debugaccess -> ROM_0:debugaccess
	wire   [9:0] mm_interconnect_1_rom_0_s1_address;         // mm_interconnect_1:ROM_0_s1_address -> ROM_0:address
	wire   [3:0] mm_interconnect_1_rom_0_s1_byteenable;      // mm_interconnect_1:ROM_0_s1_byteenable -> ROM_0:byteenable
	wire         mm_interconnect_1_rom_0_s1_write;           // mm_interconnect_1:ROM_0_s1_write -> ROM_0:write
	wire  [31:0] mm_interconnect_1_rom_0_s1_writedata;       // mm_interconnect_1:ROM_0_s1_writedata -> ROM_0:writedata
	wire         mm_interconnect_1_rom_0_s1_clken;           // mm_interconnect_1:ROM_0_s1_clken -> ROM_0:clken
	wire         irq_mapper_receiver0_irq;                   // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                   // buttons_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_0_irq_irq;                              // irq_mapper:sender_irq -> CPU_0:irq
	wire         rst_controller_reset_out_reset;             // rst_controller:reset_out -> [CPU_0:reset_n, RAM_0:reset, ROM_0:reset, buttons_0:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:CPU_0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, segm_min_0:reset_n, segm_ms_0:reset_n, segm_s_0:reset_n, switches_0:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;         // rst_controller:reset_req -> [RAM_0:reset_req, ROM_0:reset_req, rst_translator:reset_req_in]

	platform_CPU_0 cpu_0 (
		.clk           (clk_clk),                              //                       clk.clk
		.reset_n       (~rst_controller_reset_out_reset),      //                     reset.reset_n
		.d_address     (cpu_0_data_master_address),            //               data_master.address
		.d_byteenable  (cpu_0_data_master_byteenable),         //                          .byteenable
		.d_read        (cpu_0_data_master_read),               //                          .read
		.d_readdata    (cpu_0_data_master_readdata),           //                          .readdata
		.d_waitrequest (cpu_0_data_master_waitrequest),        //                          .waitrequest
		.d_write       (cpu_0_data_master_write),              //                          .write
		.d_writedata   (cpu_0_data_master_writedata),          //                          .writedata
		.i_address     (cpu_0_instruction_master_address),     //        instruction_master.address
		.i_read        (cpu_0_instruction_master_read),        //                          .read
		.i_readdata    (cpu_0_instruction_master_readdata),    //                          .readdata
		.i_waitrequest (cpu_0_instruction_master_waitrequest), //                          .waitrequest
		.irq           (cpu_0_irq_irq),                        //                       irq.irq
		.dummy_ci_port ()                                      // custom_instruction_master.readra
	);

	platform_RAM_0 ram_0 (
		.clk        (clk_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_ram_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze     (1'b0)                                   // (terminated)
	);

	platform_ROM_0 rom_0 (
		.clk         (clk_clk),                                //   clk1.clk
		.address     (mm_interconnect_1_rom_0_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_1_rom_0_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_1_rom_0_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_1_rom_0_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_1_rom_0_s1_write),       //       .write
		.readdata    (mm_interconnect_1_rom_0_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_1_rom_0_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_1_rom_0_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	platform_buttons_0 buttons_0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_buttons_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buttons_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buttons_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buttons_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buttons_0_s1_readdata),   //                    .readdata
		.in_port    (pio_0_external_connection_export),          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                   //                 irq.irq
	);

	platform_segm_min_0 segm_min_0 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_segm_min_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segm_min_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segm_min_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segm_min_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segm_min_0_s1_readdata),   //                    .readdata
		.out_port   (id7segm_min_0_external_connection_export)    // external_connection.export
	);

	platform_segm_min_0 segm_ms_0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_segm_ms_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segm_ms_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segm_ms_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segm_ms_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segm_ms_0_s1_readdata),   //                    .readdata
		.out_port   (id7segm_ms_0_external_connection_export)    // external_connection.export
	);

	platform_segm_min_0 segm_s_0 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segm_s_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segm_s_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segm_s_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segm_s_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segm_s_0_s1_readdata),   //                    .readdata
		.out_port   (id7segm_s_0_external_connection_export)    // external_connection.export
	);

	platform_switches_0 switches_0 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_switches_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_0_s1_readdata), //                    .readdata
		.in_port  (switches_0_external_connection_export)     // external_connection.export
	);

	platform_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	platform_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                           (clk_clk),                                    //                         clk_0_clk.clk
		.CPU_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),             // CPU_0_reset_reset_bridge_in_reset.reset
		.CPU_0_data_master_address               (cpu_0_data_master_address),                  //                 CPU_0_data_master.address
		.CPU_0_data_master_waitrequest           (cpu_0_data_master_waitrequest),              //                                  .waitrequest
		.CPU_0_data_master_byteenable            (cpu_0_data_master_byteenable),               //                                  .byteenable
		.CPU_0_data_master_read                  (cpu_0_data_master_read),                     //                                  .read
		.CPU_0_data_master_readdata              (cpu_0_data_master_readdata),                 //                                  .readdata
		.CPU_0_data_master_write                 (cpu_0_data_master_write),                    //                                  .write
		.CPU_0_data_master_writedata             (cpu_0_data_master_writedata),                //                                  .writedata
		.buttons_0_s1_address                    (mm_interconnect_0_buttons_0_s1_address),     //                      buttons_0_s1.address
		.buttons_0_s1_write                      (mm_interconnect_0_buttons_0_s1_write),       //                                  .write
		.buttons_0_s1_readdata                   (mm_interconnect_0_buttons_0_s1_readdata),    //                                  .readdata
		.buttons_0_s1_writedata                  (mm_interconnect_0_buttons_0_s1_writedata),   //                                  .writedata
		.buttons_0_s1_chipselect                 (mm_interconnect_0_buttons_0_s1_chipselect),  //                                  .chipselect
		.RAM_0_s1_address                        (mm_interconnect_0_ram_0_s1_address),         //                          RAM_0_s1.address
		.RAM_0_s1_write                          (mm_interconnect_0_ram_0_s1_write),           //                                  .write
		.RAM_0_s1_readdata                       (mm_interconnect_0_ram_0_s1_readdata),        //                                  .readdata
		.RAM_0_s1_writedata                      (mm_interconnect_0_ram_0_s1_writedata),       //                                  .writedata
		.RAM_0_s1_byteenable                     (mm_interconnect_0_ram_0_s1_byteenable),      //                                  .byteenable
		.RAM_0_s1_chipselect                     (mm_interconnect_0_ram_0_s1_chipselect),      //                                  .chipselect
		.RAM_0_s1_clken                          (mm_interconnect_0_ram_0_s1_clken),           //                                  .clken
		.segm_min_0_s1_address                   (mm_interconnect_0_segm_min_0_s1_address),    //                     segm_min_0_s1.address
		.segm_min_0_s1_write                     (mm_interconnect_0_segm_min_0_s1_write),      //                                  .write
		.segm_min_0_s1_readdata                  (mm_interconnect_0_segm_min_0_s1_readdata),   //                                  .readdata
		.segm_min_0_s1_writedata                 (mm_interconnect_0_segm_min_0_s1_writedata),  //                                  .writedata
		.segm_min_0_s1_chipselect                (mm_interconnect_0_segm_min_0_s1_chipselect), //                                  .chipselect
		.segm_ms_0_s1_address                    (mm_interconnect_0_segm_ms_0_s1_address),     //                      segm_ms_0_s1.address
		.segm_ms_0_s1_write                      (mm_interconnect_0_segm_ms_0_s1_write),       //                                  .write
		.segm_ms_0_s1_readdata                   (mm_interconnect_0_segm_ms_0_s1_readdata),    //                                  .readdata
		.segm_ms_0_s1_writedata                  (mm_interconnect_0_segm_ms_0_s1_writedata),   //                                  .writedata
		.segm_ms_0_s1_chipselect                 (mm_interconnect_0_segm_ms_0_s1_chipselect),  //                                  .chipselect
		.segm_s_0_s1_address                     (mm_interconnect_0_segm_s_0_s1_address),      //                       segm_s_0_s1.address
		.segm_s_0_s1_write                       (mm_interconnect_0_segm_s_0_s1_write),        //                                  .write
		.segm_s_0_s1_readdata                    (mm_interconnect_0_segm_s_0_s1_readdata),     //                                  .readdata
		.segm_s_0_s1_writedata                   (mm_interconnect_0_segm_s_0_s1_writedata),    //                                  .writedata
		.segm_s_0_s1_chipselect                  (mm_interconnect_0_segm_s_0_s1_chipselect),   //                                  .chipselect
		.switches_0_s1_address                   (mm_interconnect_0_switches_0_s1_address),    //                     switches_0_s1.address
		.switches_0_s1_readdata                  (mm_interconnect_0_switches_0_s1_readdata),   //                                  .readdata
		.timer_0_s1_address                      (mm_interconnect_0_timer_0_s1_address),       //                        timer_0_s1.address
		.timer_0_s1_write                        (mm_interconnect_0_timer_0_s1_write),         //                                  .write
		.timer_0_s1_readdata                     (mm_interconnect_0_timer_0_s1_readdata),      //                                  .readdata
		.timer_0_s1_writedata                    (mm_interconnect_0_timer_0_s1_writedata),     //                                  .writedata
		.timer_0_s1_chipselect                   (mm_interconnect_0_timer_0_s1_chipselect)     //                                  .chipselect
	);

	platform_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                           (clk_clk),                                //                         clk_0_clk.clk
		.CPU_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),         // CPU_0_reset_reset_bridge_in_reset.reset
		.CPU_0_instruction_master_address        (cpu_0_instruction_master_address),       //          CPU_0_instruction_master.address
		.CPU_0_instruction_master_waitrequest    (cpu_0_instruction_master_waitrequest),   //                                  .waitrequest
		.CPU_0_instruction_master_read           (cpu_0_instruction_master_read),          //                                  .read
		.CPU_0_instruction_master_readdata       (cpu_0_instruction_master_readdata),      //                                  .readdata
		.ROM_0_s1_address                        (mm_interconnect_1_rom_0_s1_address),     //                          ROM_0_s1.address
		.ROM_0_s1_write                          (mm_interconnect_1_rom_0_s1_write),       //                                  .write
		.ROM_0_s1_readdata                       (mm_interconnect_1_rom_0_s1_readdata),    //                                  .readdata
		.ROM_0_s1_writedata                      (mm_interconnect_1_rom_0_s1_writedata),   //                                  .writedata
		.ROM_0_s1_byteenable                     (mm_interconnect_1_rom_0_s1_byteenable),  //                                  .byteenable
		.ROM_0_s1_chipselect                     (mm_interconnect_1_rom_0_s1_chipselect),  //                                  .chipselect
		.ROM_0_s1_clken                          (mm_interconnect_1_rom_0_s1_clken),       //                                  .clken
		.ROM_0_s1_debugaccess                    (mm_interconnect_1_rom_0_s1_debugaccess)  //                                  .debugaccess
	);

	platform_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_0_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
